package mytypes_pkg is

     type my_array_t is array (1 to 7) of integer range 0 to 255;

end package mytypes_pkg;
--package body mytypes_pkg is
	
--end package body mytypes_pkg;
