--------------------------------------------------------------------------------
--! @file
--! @ingroup    RTL
--!
--! @brief      Top module
--! @date       2012-07-27
--! @author     morten@hih.au.dk     
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity top is
	port  (
		clk : in std_logic        -- input clock, xx MHz.
	);
end top;

architecture arch of top is

begin



end arch;

